module Interface ();
endmodule
