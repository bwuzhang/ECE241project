module Interface();
endmodule
